//========================================================================
// AbsDiff_4b_GL-test
//========================================================================

`include "ece2300/ece2300-test.v"

// ece2300-lint
`include "absdiff/AbsDiff_4b_GL.v"

module Top();

  //----------------------------------------------------------------------
  // Setup
  //----------------------------------------------------------------------

  CombinationalTestUtils t();

  //----------------------------------------------------------------------
  // Instantiate design under test
  //----------------------------------------------------------------------

  logic [3:0] in0;
  logic [3:0] in1;
  logic [3:0] diff;

  AbsDiff_4b_GL dut
  (
    .in0  (in0),
    .in1  (in1),
    .diff (diff)
  );

  //----------------------------------------------------------------------
  // Include test cases
  //----------------------------------------------------------------------

  `include "absdiff/test/AbsDiff_4b-test-cases.v"

endmodule

